interface simple_if;
logic a;
logic b;
endinterface