module use_if(simple_if s);
always_comb begin
    s.b = s.a;
end
endmodule
